// ============================================================================
// mp64_mul_asic.v — ASIC Multiplier Stub
// ============================================================================
// Replace body with DesignWare DW02_mult or foundry multiplier macro.
// Port interface identical to rtl/prim/mp64_mul.v.
//

module mp64_mul #(
    parameter LATENCY = 4
)(
    input  wire         clk,
    input  wire         rst,
    input  wire         start,
    input  wire         is_signed,
    input  wire [63:0]  a,
    input  wire [63:0]  b,
    output wire [127:0] result,
    output wire         done,
    output wire         busy
);

    // STUB — behavioural fallback (replace with DW02_mult pipeline)
    reg [127:0] pipe_data [0:LATENCY-1];
    reg [LATENCY-1:0] pipe_valid;

    wire [127:0] product = is_signed
        ? $signed(a) * $signed(b)
        : a * b;

    integer i;
    always @(posedge clk) begin
        if (rst) begin
            pipe_valid <= {LATENCY{1'b0}};
            for (i = 0; i < LATENCY; i = i + 1)
                pipe_data[i] <= 128'd0;
        end else begin
            pipe_valid[0] <= start;
            pipe_data[0]  <= start ? product : pipe_data[0];
            for (i = 1; i < LATENCY; i = i + 1) begin
                pipe_valid[i] <= pipe_valid[i-1];
                pipe_data[i]  <= pipe_data[i-1];
            end
        end
    end

    assign result = pipe_data[LATENCY-1];
    assign done   = pipe_valid[LATENCY-1];
    assign busy   = start | (|pipe_valid);

endmodule
