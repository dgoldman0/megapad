// ============================================================================
// tb_field_alu.v — Field ALU Accelerator Unit Tests
// ============================================================================
//
// Tests:
//   1. FADD: (3 + 5) mod p = 8
//   2. FSUB: (5 - 3) mod p = 2
//   3. FSUB wraparound: (3 - 5) mod p = p - 2
//   4. FMUL: (7 × 11) mod p = 77
//   5. FSQR: 9² mod p = 81
//   6. FINV: inv(2) × 2 mod p = 1 (verify via readback)
//   7. MUL_RAW: 0xFF...FF × 2 → 512-bit result with overflow
//   8. X25519: scalar = 1 (clamped), base point 9 → known result
//   9. Status transitions: idle → busy → done
//  10. FPOW: 2^10 mod p = 1024
//

`timescale 1ns / 1ps
`include "mp64_defs.vh"

module tb_field_alu;

    reg clk, rst_n;
    initial clk = 0;
    always #5 clk = ~clk;  // 100 MHz

    integer pass_count = 0;
    integer fail_count = 0;
    integer test_num   = 0;

    // DUT signals
    reg         req;
    reg  [5:0]  addr;
    reg  [63:0] wdata;
    reg         wen;
    wire [63:0] rdata;
    wire        ack;

    mp64_field_alu u_dut (
        .clk(clk), .rst_n(rst_n),
        .req(req), .addr(addr), .wdata(wdata), .wen(wen),
        .rdata(rdata), .ack(ack)
    );

    // ========================================================================
    // Helper tasks
    // ========================================================================

    task write64(input [5:0] a, input [63:0] d);
        begin
            @(posedge clk);
            req <= 1; addr <= a; wdata <= d; wen <= 1;
            @(posedge clk);
            req <= 0; wen <= 0;
        end
    endtask

    task read64(input [5:0] a, output [63:0] d);
        begin
            @(posedge clk);
            req <= 1; addr <= a; wdata <= 0; wen <= 0;
            @(posedge clk);
            req <= 0;
            @(posedge clk);  // wait for registered rdata to settle
            d = rdata;
        end
    endtask

    // Write 256-bit operand A (4 × 64-bit LE words)
    task write_operand_a(input [255:0] val);
        begin
            write64(6'h00, val[ 63:  0]);
            write64(6'h08, val[127: 64]);
            write64(6'h10, val[191:128]);
            write64(6'h18, val[255:192]);
        end
    endtask

    // Write 256-bit operand B
    task write_operand_b(input [255:0] val);
        begin
            write64(6'h20, val[ 63:  0]);
            write64(6'h28, val[127: 64]);
            write64(6'h30, val[191:128]);
            write64(6'h38, val[255:192]);
        end
    endtask

    // Issue CMD: mode in bits [4:1], go in bit [0], result_sel in bit [5]
    task issue_cmd(input [3:0] mode, input go, input result_sel);
        begin
            write64(6'h3F, {58'd0, result_sel, mode, go});
        end
    endtask

    // Wait for done (polls STATUS until done bit = 1)
    task wait_done;
        reg [63:0] st;
        integer timeout;
        begin
            timeout = 0;
            st = 0;
            while (!st[1] && timeout < 200000) begin
                read64(6'h00, st);
                timeout = timeout + 1;
            end
            if (timeout >= 200000) begin
                $display("  TIMEOUT waiting for done!");
                fail_count = fail_count + 1;
            end
        end
    endtask

    // Read 256-bit result (LO or HI depending on result_sel)
    task read_result(output [255:0] val);
        reg [63:0] w0, w1, w2, w3;
        begin
            read64(6'h08, w0);
            read64(6'h10, w1);
            read64(6'h18, w2);
            read64(6'h20, w3);
            val = {w3, w2, w1, w0};
        end
    endtask

    // Check helper
    task check(input [255:0] got, input [255:0] expected, input [8*40-1:0] name);
        begin
            test_num = test_num + 1;
            if (got === expected) begin
                $display("  [PASS] Test %0d: %0s", test_num, name);
                pass_count = pass_count + 1;
            end else begin
                $display("  [FAIL] Test %0d: %0s", test_num, name);
                $display("         expected: %064h", expected);
                $display("              got: %064h", got);
                fail_count = fail_count + 1;
            end
        end
    endtask

    // ========================================================================
    // Test sequence
    // ========================================================================
    reg [255:0] result;
    reg [63:0]  status;

    localparam [255:0] PRIME = 256'h7FFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFFF_FFFFFFED;

    initial begin
        $dumpfile("tb_field_alu.vcd");
        $dumpvars(0, tb_field_alu);

        req <= 0; addr <= 0; wdata <= 0; wen <= 0;
        rst_n = 0;
        #20;
        rst_n = 1;
        #10;

        $display("=== Field ALU Tests ===");

        // --- Test 1: FADD (3 + 5) = 8 ---
        write_operand_a(256'd3);
        write_operand_b(256'd5);
        issue_cmd(4'd1, 1'b1, 1'b0);  // mode=FADD, go
        wait_done;
        read_result(result);
        check(result, 256'd8, "FADD(3,5)=8");

        // --- Test 2: FSUB (5 - 3) = 2 ---
        write_operand_a(256'd5);
        write_operand_b(256'd3);
        issue_cmd(4'd2, 1'b1, 1'b0);  // FSUB
        wait_done;
        read_result(result);
        check(result, 256'd2, "FSUB(5,3)=2");

        // --- Test 3: FSUB wraparound (3 - 5) mod p = p - 2 ---
        write_operand_a(256'd3);
        write_operand_b(256'd5);
        issue_cmd(4'd2, 1'b1, 1'b0);
        wait_done;
        read_result(result);
        check(result, PRIME - 256'd2, "FSUB(3,5)=p-2");

        // --- Test 4: FMUL (7 × 11) = 77 ---
        write_operand_a(256'd7);
        write_operand_b(256'd11);
        issue_cmd(4'd3, 1'b1, 1'b0);  // FMUL
        wait_done;
        read_result(result);
        check(result, 256'd77, "FMUL(7,11)=77");

        // --- Test 5: FSQR (9²) = 81 ---
        write_operand_a(256'd9);
        issue_cmd(4'd4, 1'b1, 1'b0);  // FSQR
        wait_done;
        read_result(result);
        check(result, 256'd81, "FSQR(9)=81");

        // --- Test 6: FINV — compute 2⁻¹ mod p ---
        // p = 2²⁵⁵ − 19, so 2⁻¹ = (p+1)/2
        write_operand_a(256'd2);
        issue_cmd(4'd5, 1'b1, 1'b0);  // FINV
        wait_done;
        read_result(result);
        check(result, (PRIME + 256'd1) >> 1, "FINV(2)=(p+1)/2");

        // --- Test 7: MUL_RAW — small values, verify low half ---
        write_operand_a(256'd100);
        write_operand_b(256'd200);
        issue_cmd(4'd7, 1'b1, 1'b0);  // MUL_RAW
        wait_done;
        read_result(result);  // reads LO (result_sel=0)
        check(result, 256'd20000, "MUL_RAW(100,200) LO=20000");

        // Read HI half (should be 0 for small operands)
        issue_cmd(4'd0, 1'b0, 1'b1);  // set result_sel=1, no go
        @(posedge clk); @(posedge clk);
        read_result(result);
        check(result, 256'd0, "MUL_RAW(100,200) HI=0");

        // --- Test 8: Status — verify idle→busy→done ---
        // Already done, just verify status reads done
        issue_cmd(4'd0, 1'b0, 1'b0);  // reset result_sel
        @(posedge clk);
        read64(6'h00, status);
        check({192'd0, status}, {192'd0, 62'd0, 2'b10}, "STATUS=done(2)");

        // --- Test 9: FPOW — 2^10 mod p = 1024 ---
        write_operand_a(256'd2);
        write_operand_b(256'd10);
        issue_cmd(4'd6, 1'b1, 1'b0);  // FPOW
        wait_done;
        read_result(result);
        check(result, 256'd1024, "FPOW(2,10)=1024");

        // --- Test 10: FMUL identity — a × 1 = a (a < p) ---
        write_operand_a(256'h1EADBEEF_CAFEBABE_12345678_9ABCDEF0_DEADBEEF_CAFEBABE_12345678_9ABCDEF0);
        write_operand_b(256'd1);
        issue_cmd(4'd3, 1'b1, 1'b0);  // FMUL
        wait_done;
        read_result(result);
        check(result, 256'h1EADBEEF_CAFEBABE_12345678_9ABCDEF0_DEADBEEF_CAFEBABE_12345678_9ABCDEF0,
              "FMUL(x,1)=x");

        // ================================================================
        $display("");
        $display("=== Results: %0d passed, %0d failed ===", pass_count, fail_count);
        if (fail_count == 0)
            $display("ALL TESTS PASSED");
        else
            $display("SOME TESTS FAILED");
        $finish;
    end

endmodule
